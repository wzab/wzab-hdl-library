library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

package genlfsr_pkg is

  type T_LFSR_TAPS is array (natural range <>) of integer;

end genlfsr_pkg;
